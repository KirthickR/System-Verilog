interface intf;
  logic d;
  logic clk;
  logic rst;
  logic q;
  logic qbar;
endinterface
